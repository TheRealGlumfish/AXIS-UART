../../rtl/uart.vhd